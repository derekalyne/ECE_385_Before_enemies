module intial_enemy_dug(input               Clk,
								input [23:0]        update_dug_state[31:0],
								output [23:0]       dug_state[31:0]);
		
endmodule 